module ROM(Addr,Dout);
    input [9:0] Addr;
    output reg [31:0] Dout;
    always@(Addr)begin
        case(Addr)
            10'b0000000000 :Dout=32'h00100493;
            10'b0000000001 :Dout=32'h0100006f;
            10'b0000000010 :Dout=32'h00100493;
            10'b0000000011 :Dout=32'h00200913;
            10'b0000000100 :Dout=32'h00300993;
            10'b0000000101 :Dout=32'h0100006f;
            10'b0000000110 :Dout=32'h00100493;
            10'b0000000111 :Dout=32'h00200913;
            10'b0000001000 :Dout=32'h00300993;
            10'b0000001001 :Dout=32'h0100006f;
            10'b0000001010 :Dout=32'h00100493;
            10'b0000001011 :Dout=32'h00200913;
            10'b0000001100 :Dout=32'h00300993;
            10'b0000001101 :Dout=32'h0100006f;
            10'b0000001110 :Dout=32'h00100493;
            10'b0000001111 :Dout=32'h00200913;
            10'b0000010000 :Dout=32'h00300993;
            10'b0000010001 :Dout=32'h3a0000ef;
            10'b0000010010 :Dout=32'h00100413;
            10'b0000010011 :Dout=32'h00100493;
            10'b0000010100 :Dout=32'h01f49493;
            10'b0000010101 :Dout=32'h00900533;
            10'b0000010110 :Dout=32'h02200893;
            10'b0000010111 :Dout=32'h00000073;
            10'b0000011000 :Dout=32'h0024d493;
            10'b0000011001 :Dout=32'h00048463;
            10'b0000011010 :Dout=32'hfedff06f;
            10'b0000011011 :Dout=32'h00900533;
            10'b0000011100 :Dout=32'h02200893;
            10'b0000011101 :Dout=32'h00000073;
            10'b0000011110 :Dout=32'h00100493;
            10'b0000011111 :Dout=32'h00249493;
            10'b0000100000 :Dout=32'h00900533;
            10'b0000100001 :Dout=32'h02200893;
            10'b0000100010 :Dout=32'h00000073;
            10'b0000100011 :Dout=32'h00048463;
            10'b0000100100 :Dout=32'hfedff06f;
            10'b0000100101 :Dout=32'h00100493;
            10'b0000100110 :Dout=32'h01f49493;
            10'b0000100111 :Dout=32'h00900533;
            10'b0000101000 :Dout=32'h02200893;
            10'b0000101001 :Dout=32'h00000073;
            10'b0000101010 :Dout=32'h4034d493;
            10'b0000101011 :Dout=32'h00900533;
            10'b0000101100 :Dout=32'h02200893;
            10'b0000101101 :Dout=32'h00000073;
            10'b0000101110 :Dout=32'h4044d493;
            10'b0000101111 :Dout=32'h00900533;
            10'b0000110000 :Dout=32'h02200893;
            10'b0000110001 :Dout=32'h00000073;
            10'b0000110010 :Dout=32'h4044d493;
            10'b0000110011 :Dout=32'h00900533;
            10'b0000110100 :Dout=32'h02200893;
            10'b0000110101 :Dout=32'h00000073;
            10'b0000110110 :Dout=32'h4044d493;
            10'b0000110111 :Dout=32'h00900533;
            10'b0000111000 :Dout=32'h02200893;
            10'b0000111001 :Dout=32'h00000073;
            10'b0000111010 :Dout=32'h4044d493;
            10'b0000111011 :Dout=32'h00900533;
            10'b0000111100 :Dout=32'h02200893;
            10'b0000111101 :Dout=32'h00000073;
            10'b0000111110 :Dout=32'h4044d493;
            10'b0000111111 :Dout=32'h00900533;
            10'b0001000000 :Dout=32'h02200893;
            10'b0001000001 :Dout=32'h00000073;
            10'b0001000010 :Dout=32'h4044d493;
            10'b0001000011 :Dout=32'h00900533;
            10'b0001000100 :Dout=32'h02200893;
            10'b0001000101 :Dout=32'h00000073;
            10'b0001000110 :Dout=32'h4044d493;
            10'b0001000111 :Dout=32'h00900533;
            10'b0001001000 :Dout=32'h02200893;
            10'b0001001001 :Dout=32'h00000073;
            10'b0001001010 :Dout=32'h00100413;
            10'b0001001011 :Dout=32'h01f41993;
            10'b0001001100 :Dout=32'h41f9d993;
            10'b0001001101 :Dout=32'h00000433;
            10'b0001001110 :Dout=32'h00c00913;
            10'b0001001111 :Dout=32'h00300b13;
            10'b0001010000 :Dout=32'h00140413;
            10'b0001010001 :Dout=32'h00f47413;
            10'b0001010010 :Dout=32'h00800293;
            10'b0001010011 :Dout=32'h00100313;
            10'b0001010100 :Dout=32'h00499993;
            10'b0001010101 :Dout=32'h0089e9b3;
            10'b0001010110 :Dout=32'h01300533;
            10'b0001010111 :Dout=32'h02200893;
            10'b0001011000 :Dout=32'h00000073;
            10'b0001011001 :Dout=32'h406282b3;
            10'b0001011010 :Dout=32'hfe0294e3;
            10'b0001011011 :Dout=32'h00140413;
            10'b0001011100 :Dout=32'h00f00f93;
            10'b0001011101 :Dout=32'h01f47433;
            10'b0001011110 :Dout=32'h01c41413;
            10'b0001011111 :Dout=32'h00800293;
            10'b0001100000 :Dout=32'h00100313;
            10'b0001100001 :Dout=32'h0049d993;
            10'b0001100010 :Dout=32'h0089e9b3;
            10'b0001100011 :Dout=32'h01300533;
            10'b0001100100 :Dout=32'h02200893;
            10'b0001100101 :Dout=32'h00000073;
            10'b0001100110 :Dout=32'h406282b3;
            10'b0001100111 :Dout=32'hfe0294e3;
            10'b0001101000 :Dout=32'h01c45413;
            10'b0001101001 :Dout=32'h406b0b33;
            10'b0001101010 :Dout=32'h000b0463;
            10'b0001101011 :Dout=32'hf95ff06f;
            10'b0001101100 :Dout=32'h000002b3;
            10'b0001101101 :Dout=32'hfff2c293;
            10'b0001101110 :Dout=32'h00829293;
            10'b0001101111 :Dout=32'h0ff2e293;
            10'b0001110000 :Dout=32'h00500533;
            10'b0001110001 :Dout=32'h02200893;
            10'b0001110010 :Dout=32'h00000073;
            10'b0001110011 :Dout=32'hfff00413;
            10'b0001110100 :Dout=32'h00000493;
            10'b0001110101 :Dout=32'h0084a023;
            10'b0001110110 :Dout=32'h00140413;
            10'b0001110111 :Dout=32'h00448493;
            10'b0001111000 :Dout=32'h0084a023;
            10'b0001111001 :Dout=32'h00140413;
            10'b0001111010 :Dout=32'h00448493;
            10'b0001111011 :Dout=32'h0084a023;
            10'b0001111100 :Dout=32'h00140413;
            10'b0001111101 :Dout=32'h00448493;
            10'b0001111110 :Dout=32'h0084a023;
            10'b0001111111 :Dout=32'h00140413;
            10'b0010000000 :Dout=32'h00448493;
            10'b0010000001 :Dout=32'h0084a023;
            10'b0010000010 :Dout=32'h00140413;
            10'b0010000011 :Dout=32'h00448493;
            10'b0010000100 :Dout=32'h0084a023;
            10'b0010000101 :Dout=32'h00140413;
            10'b0010000110 :Dout=32'h00448493;
            10'b0010000111 :Dout=32'h0084a023;
            10'b0010001000 :Dout=32'h00140413;
            10'b0010001001 :Dout=32'h00448493;
            10'b0010001010 :Dout=32'h0084a023;
            10'b0010001011 :Dout=32'h00140413;
            10'b0010001100 :Dout=32'h00448493;
            10'b0010001101 :Dout=32'h0084a023;
            10'b0010001110 :Dout=32'h00140413;
            10'b0010001111 :Dout=32'h00448493;
            10'b0010010000 :Dout=32'h0084a023;
            10'b0010010001 :Dout=32'h00140413;
            10'b0010010010 :Dout=32'h00448493;
            10'b0010010011 :Dout=32'h0084a023;
            10'b0010010100 :Dout=32'h00140413;
            10'b0010010101 :Dout=32'h00448493;
            10'b0010010110 :Dout=32'h0084a023;
            10'b0010010111 :Dout=32'h00140413;
            10'b0010011000 :Dout=32'h00448493;
            10'b0010011001 :Dout=32'h0084a023;
            10'b0010011010 :Dout=32'h00140413;
            10'b0010011011 :Dout=32'h00448493;
            10'b0010011100 :Dout=32'h0084a023;
            10'b0010011101 :Dout=32'h00140413;
            10'b0010011110 :Dout=32'h00448493;
            10'b0010011111 :Dout=32'h0084a023;
            10'b0010100000 :Dout=32'h00140413;
            10'b0010100001 :Dout=32'h00448493;
            10'b0010100010 :Dout=32'h0084a023;
            10'b0010100011 :Dout=32'h00140413;
            10'b0010100100 :Dout=32'h00448493;
            10'b0010100101 :Dout=32'h00140413;
            10'b0010100110 :Dout=32'h00000433;
            10'b0010100111 :Dout=32'h03c00493;
            10'b0010101000 :Dout=32'h00042983;
            10'b0010101001 :Dout=32'h0004aa03;
            10'b0010101010 :Dout=32'h0149a2b3;
            10'b0010101011 :Dout=32'h00028663;
            10'b0010101100 :Dout=32'h0134a023;
            10'b0010101101 :Dout=32'h01442023;
            10'b0010101110 :Dout=32'hffc48493;
            10'b0010101111 :Dout=32'hfe9412e3;
            10'b0010110000 :Dout=32'h00800533;
            10'b0010110001 :Dout=32'h02200893;
            10'b0010110010 :Dout=32'h00000073;
            10'b0010110011 :Dout=32'h00440413;
            10'b0010110100 :Dout=32'h03c00493;
            10'b0010110101 :Dout=32'hfc9416e3;
            10'b0010110110 :Dout=32'h03200893;
            10'b0010110111 :Dout=32'h00000073;
            10'b0010111000 :Dout=32'h00100293;
            10'b0010111001 :Dout=32'h00300313;
            10'b0010111010 :Dout=32'h00800493;
            10'b0010111011 :Dout=32'h00849493;
            10'b0010111100 :Dout=32'h07648493;
            10'b0010111101 :Dout=32'h01449493;
            10'b0010111110 :Dout=32'h00900533;
            10'b0010111111 :Dout=32'h02200893;
            10'b0011000000 :Dout=32'h00000073;
            10'b0011000001 :Dout=32'h00800e13;
            10'b0011000010 :Dout=32'h0054d4b3;
            10'b0011000011 :Dout=32'h0064d4b3;
            10'b0011000100 :Dout=32'h00900533;
            10'b0011000101 :Dout=32'h02200893;
            10'b0011000110 :Dout=32'h00000073;
            10'b0011000111 :Dout=32'hfffe0e13;
            10'b0011001000 :Dout=32'hfe0e14e3;
            10'b0011001001 :Dout=32'h00a00893;
            10'b0011001010 :Dout=32'h00000073;
            10'b0011001011 :Dout=32'hfff00293;
            10'b0011001100 :Dout=32'h00000313;
            10'b0011001101 :Dout=32'h01900413;
            10'b0011001110 :Dout=32'h00841413;
            10'b0011001111 :Dout=32'h09700493;
            10'b0011010000 :Dout=32'h00940533;
            10'b0011010001 :Dout=32'h02200893;
            10'b0011010010 :Dout=32'h00000073;
            10'b0011010011 :Dout=32'h005484b3;
            10'b0011010100 :Dout=32'h0494b313;
            10'b0011010101 :Dout=32'hfe0306e3;
            10'b0011010110 :Dout=32'h00a00893;
            10'b0011010111 :Dout=32'h00000073;
            10'b0011011000 :Dout=32'h00000313;
            10'b0011011001 :Dout=32'h02000e13;
            10'b0011011010 :Dout=32'h00000493;
            10'b0011011011 :Dout=32'h00100913;
            10'b0011011100 :Dout=32'h00930023;
            10'b0011011101 :Dout=32'h00900533;
            10'b0011011110 :Dout=32'h02200893;
            10'b0011011111 :Dout=32'h00000073;
            10'b0011100000 :Dout=32'h012484b3;
            10'b0011100001 :Dout=32'h00130313;
            10'b0011100010 :Dout=32'hfffe0e13;
            10'b0011100011 :Dout=32'hfe0e12e3;
            10'b0011100100 :Dout=32'h00800e13;
            10'b0011100101 :Dout=32'h00000313;
            10'b0011100110 :Dout=32'h00032483;
            10'b0011100111 :Dout=32'h00900533;
            10'b0011101000 :Dout=32'h02200893;
            10'b0011101001 :Dout=32'h00000073;
            10'b0011101010 :Dout=32'h00430313;
            10'b0011101011 :Dout=32'hfffe0e13;
            10'b0011101100 :Dout=32'hfe0e14e3;
            10'b0011101101 :Dout=32'h00a00893;
            10'b0011101110 :Dout=32'h00000073;
            10'b0011101111 :Dout=32'hff100493;
            10'b0011110000 :Dout=32'h00900533;
            10'b0011110001 :Dout=32'h02200893;
            10'b0011110010 :Dout=32'h00000073;
            10'b0011110011 :Dout=32'h00148493;
            10'b0011110100 :Dout=32'hfe04c8e3;
            10'b0011110101 :Dout=32'h00a00893;
            10'b0011110110 :Dout=32'h00000073;
            10'b0011110111 :Dout=32'h00a00893;
            10'b0011111000 :Dout=32'h00000073;
            10'b0011111001 :Dout=32'h00000413;
            10'b0011111010 :Dout=32'h00140413;
            10'b0011111011 :Dout=32'h00800533;
            10'b0011111100 :Dout=32'h02200893;
            10'b0011111101 :Dout=32'h00000073;
            10'b0011111110 :Dout=32'h00240413;
            10'b0011111111 :Dout=32'h00800533;
            10'b0100000000 :Dout=32'h02200893;
            10'b0100000001 :Dout=32'h00000073;
            10'b0100000010 :Dout=32'h00340413;
            10'b0100000011 :Dout=32'h00800533;
            10'b0100000100 :Dout=32'h02200893;
            10'b0100000101 :Dout=32'h00000073;
            10'b0100000110 :Dout=32'h00440413;
            10'b0100000111 :Dout=32'h00800533;
            10'b0100001000 :Dout=32'h02200893;
            10'b0100001001 :Dout=32'h00000073;
            10'b0100001010 :Dout=32'h00540413;
            10'b0100001011 :Dout=32'h00800533;
            10'b0100001100 :Dout=32'h02200893;
            10'b0100001101 :Dout=32'h00000073;
            10'b0100001110 :Dout=32'h00640413;
            10'b0100001111 :Dout=32'h00800533;
            10'b0100010000 :Dout=32'h02200893;
            10'b0100010001 :Dout=32'h00000073;
            10'b0100010010 :Dout=32'h00740413;
            10'b0100010011 :Dout=32'h00800533;
            10'b0100010100 :Dout=32'h02200893;
            10'b0100010101 :Dout=32'h00000073;
            10'b0100010110 :Dout=32'h00840413;
            10'b0100010111 :Dout=32'h00800533;
            10'b0100011000 :Dout=32'h02200893;
            10'b0100011001 :Dout=32'h02200893;
            10'b0100011010 :Dout=32'h00000073;
            10'b0100011011 :Dout=32'h00008067;
            default: Dout=0;
        endcase
    end
endmodule